library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.all;

entity maths is
port (clk : in std_logic;
      o_sel	: in std_logic;
        data_i : in std_logic_vector(9 downto 0);
        data_o : out std_logic_vector(9 downto 0);
		ir_in	: in std_logic_vector(9 downto 0);
		red_in	: in std_logic_vector(9 downto 0);
		  set_mode: out std_logic;
		  sw_in : in std_logic
     );
end maths;
--GOOD
architecture Behavioral of maths is

--Declaration of type and signal of a 256 element RAM
--with each element being 8 bit wide.
signal sclk : std_logic := '0';
signal red : integer := 0;
signal ir : integer := 0;
signal temp : std_logic_vector (9 downto 0) := "0000000000";
signal temp2 : std_logic_vector (9 downto 0) := "0000000000";
signal four : std_logic_vector (9 downto 0) := "0000000100";
signal red_int : std_logic_vector(9 downto 0);
signal ir_int :  std_logic_vector(9 downto 0);
signal switch : std_logic := '0';
signal index : integer := 0;
signal last_sat : std_logic_vector(9 downto 0) := "0001100011";
signal avg_sat : std_logic_vector(9 downto 0) := "0000000000";
signal cur_sat : std_logic_vector(9 downto 0) := "0000000000";
signal sum_sat : std_logic_vector(9 downto 0) := "0000000000";
type ram_sat is array (0 to 2303) of std_logic_vector(7 downto 0);
type ram_ir is array (0 to 47) of std_logic_vector (11 downto 0);
signal sat: ram_sat := (X"63",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"43",X"2F",X"29",X"25",X"22",X"20",X"1F",X"1E",X"1D",X"1C",X"1C",X"1B",X"1B",X"1A",X"1A",X"19",X"19",X"19",X"18",X"18",X"18",X"18",X"17",X"17",X"17",X"17",X"17",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"14",X"14",X"14",X"63",X"5D",X"43",X"39",X"34",X"30",X"2E",X"2C",X"2A",X"29",X"28",X"27",X"26",X"25",X"25",X"24",X"24",X"23",X"23",X"22",X"22",X"22",X"21",X"21",X"21",X"20",X"20",X"20",X"20",X"1F",X"1F",X"1F",X"1F",X"1F",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"63",X"63",X"4E",X"43",X"3C",X"38",X"35",X"33",X"31",X"30",X"2F",X"2D",X"2C",X"2C",X"2B",X"2A",X"2A",X"29",X"29",X"28",X"28",X"27",X"27",X"26",X"26",X"26",X"26",X"25",X"25",X"25",X"24",X"24",X"24",X"24",X"24",X"23",X"23",X"23",X"23",X"23",X"23",X"22",X"22",X"22",X"22",X"22",X"22",X"21",X"63",X"63",X"56",X"49",X"43",X"3E",X"3B",X"38",X"36",X"35",X"33",X"32",X"31",X"30",X"2F",X"2F",X"2E",X"2D",X"2D",X"2C",X"2C",X"2B",X"2B",X"2A",X"2A",X"2A",X"29",X"29",X"29",X"28",X"28",X"28",X"28",X"27",X"27",X"27",X"27",X"27",X"26",X"26",X"26",X"26",X"26",X"26",X"25",X"25",X"25",X"25",X"63",X"63",X"5C",X"4F",X"47",X"43",X"3F",X"3C",X"3A",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"31",X"30",X"2F",X"2F",X"2E",X"2E",X"2E",X"2D",X"2D",X"2C",X"2C",X"2C",X"2B",X"2B",X"2B",X"2B",X"2A",X"2A",X"2A",X"2A",X"29",X"29",X"29",X"29",X"29",X"28",X"28",X"28",X"28",X"28",X"28",X"63",X"63",X"61",X"53",X"4B",X"46",X"43",X"40",X"3D",X"3C",X"3A",X"39",X"38",X"36",X"36",X"35",X"34",X"33",X"33",X"32",X"31",X"31",X"30",X"30",X"30",X"2F",X"2F",X"2E",X"2E",X"2E",X"2E",X"2D",X"2D",X"2D",X"2C",X"2C",X"2C",X"2C",X"2B",X"2B",X"2B",X"2B",X"2B",X"2A",X"2A",X"2A",X"2A",X"2A",X"63",X"63",X"63",X"57",X"4F",X"49",X"45",X"43",X"40",X"3E",X"3D",X"3B",X"3A",X"39",X"38",X"37",X"36",X"35",X"35",X"34",X"34",X"33",X"33",X"32",X"32",X"31",X"31",X"31",X"30",X"30",X"30",X"2F",X"2F",X"2F",X"2E",X"2E",X"2E",X"2E",X"2D",X"2D",X"2D",X"2D",X"2D",X"2C",X"2C",X"2C",X"2C",X"2C",X"63",X"63",X"63",X"5A",X"51",X"4C",X"48",X"45",X"43",X"41",X"3F",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"37",X"37",X"36",X"36",X"35",X"34",X"34",X"34",X"33",X"33",X"32",X"32",X"32",X"31",X"31",X"31",X"30",X"30",X"30",X"30",X"2F",X"2F",X"2F",X"2F",X"2E",X"2E",X"2E",X"2E",X"2E",X"2D",X"2D",X"63",X"63",X"63",X"5D",X"54",X"4E",X"4A",X"47",X"45",X"43",X"41",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"38",X"37",X"37",X"36",X"36",X"35",X"35",X"34",X"34",X"34",X"33",X"33",X"32",X"32",X"32",X"32",X"31",X"31",X"31",X"31",X"30",X"30",X"30",X"30",X"2F",X"2F",X"2F",X"2F",X"2F",X"63",X"63",X"63",X"5F",X"56",X"50",X"4C",X"49",X"46",X"44",X"43",X"41",X"40",X"3E",X"3D",X"3C",X"3C",X"3B",X"3A",X"39",X"39",X"38",X"38",X"37",X"37",X"36",X"36",X"35",X"35",X"35",X"34",X"34",X"34",X"33",X"33",X"33",X"32",X"32",X"32",X"32",X"31",X"31",X"31",X"31",X"31",X"30",X"30",X"30",X"63",X"63",X"63",X"61",X"58",X"52",X"4E",X"4B",X"48",X"46",X"44",X"43",X"41",X"40",X"3F",X"3E",X"3D",X"3C",X"3B",X"3B",X"3A",X"39",X"39",X"38",X"38",X"37",X"37",X"37",X"36",X"36",X"35",X"35",X"35",X"34",X"34",X"34",X"34",X"33",X"33",X"33",X"33",X"32",X"32",X"32",X"32",X"31",X"31",X"31",X"63",X"63",X"63",X"63",X"5A",X"54",X"50",X"4C",X"4A",X"47",X"46",X"44",X"43",X"41",X"40",X"3F",X"3E",X"3D",X"3D",X"3C",X"3B",X"3B",X"3A",X"3A",X"39",X"39",X"38",X"38",X"37",X"37",X"37",X"36",X"36",X"36",X"35",X"35",X"35",X"34",X"34",X"34",X"34",X"33",X"33",X"33",X"33",X"33",X"32",X"32",X"63",X"63",X"63",X"63",X"5C",X"56",X"51",X"4E",X"4B",X"49",X"47",X"45",X"44",X"43",X"41",X"40",X"3F",X"3F",X"3E",X"3D",X"3C",X"3C",X"3B",X"3B",X"3A",X"3A",X"39",X"39",X"38",X"38",X"38",X"37",X"37",X"37",X"36",X"36",X"36",X"35",X"35",X"35",X"35",X"34",X"34",X"34",X"34",X"33",X"33",X"33",X"63",X"63",X"63",X"63",X"5D",X"57",X"53",X"4F",X"4C",X"4A",X"48",X"46",X"45",X"44",X"43",X"41",X"41",X"40",X"3F",X"3E",X"3D",X"3D",X"3C",X"3C",X"3B",X"3B",X"3A",X"3A",X"39",X"39",X"39",X"38",X"38",X"38",X"37",X"37",X"37",X"36",X"36",X"36",X"36",X"35",X"35",X"35",X"35",X"34",X"34",X"34",X"63",X"63",X"63",X"63",X"5F",X"59",X"54",X"50",X"4E",X"4B",X"49",X"48",X"46",X"45",X"44",X"43",X"42",X"41",X"40",X"3F",X"3E",X"3E",X"3D",X"3D",X"3C",X"3C",X"3B",X"3B",X"3A",X"3A",X"39",X"39",X"39",X"38",X"38",X"38",X"37",X"37",X"37",X"37",X"36",X"36",X"36",X"36",X"35",X"35",X"35",X"35",X"63",X"63",X"63",X"63",X"60",X"5A",X"55",X"52",X"4F",X"4C",X"4A",X"49",X"47",X"46",X"45",X"43",X"43",X"42",X"41",X"40",X"3F",X"3F",X"3E",X"3E",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"38",X"38",X"38",X"37",X"37",X"37",X"37",X"36",X"36",X"36",X"36",X"36",X"63",X"63",X"63",X"63",X"62",X"5B",X"56",X"53",X"50",X"4D",X"4B",X"4A",X"48",X"47",X"45",X"44",X"43",X"43",X"42",X"41",X"40",X"40",X"3F",X"3E",X"3E",X"3D",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"38",X"38",X"38",X"38",X"37",X"37",X"37",X"37",X"37",X"36",X"63",X"63",X"63",X"63",X"63",X"5C",X"57",X"54",X"51",X"4E",X"4C",X"4B",X"49",X"48",X"46",X"45",X"44",X"43",X"43",X"42",X"41",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3D",X"3D",X"3C",X"3C",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"39",X"38",X"38",X"38",X"38",X"37",X"37",X"37",X"63",X"63",X"63",X"63",X"63",X"5D",X"58",X"55",X"52",X"4F",X"4D",X"4B",X"4A",X"48",X"47",X"46",X"45",X"44",X"43",X"43",X"42",X"41",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"39",X"38",X"38",X"38",X"38",X"63",X"63",X"63",X"63",X"63",X"5E",X"59",X"56",X"53",X"50",X"4E",X"4C",X"4B",X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"43",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3D",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"39",X"38",X"38",X"63",X"63",X"63",X"63",X"63",X"5F",X"5A",X"57",X"53",X"51",X"4F",X"4D",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"44",X"43",X"43",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"3A",X"39",X"39",X"39",X"63",X"63",X"63",X"63",X"63",X"60",X"5B",X"57",X"54",X"52",X"50",X"4E",X"4C",X"4B",X"49",X"48",X"47",X"46",X"45",X"45",X"44",X"43",X"43",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"3A",X"39",X"63",X"63",X"63",X"63",X"63",X"61",X"5C",X"58",X"55",X"53",X"50",X"4E",X"4D",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"45",X"44",X"43",X"43",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3A",X"3A",X"3A",X"63",X"63",X"63",X"63",X"63",X"62",X"5D",X"59",X"56",X"53",X"51",X"4F",X"4E",X"4C",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",X"44",X"44",X"43",X"43",X"42",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"3B",X"3A",X"63",X"63",X"63",X"63",X"63",X"63",X"5E",X"5A",X"57",X"54",X"52",X"50",X"4E",X"4D",X"4B",X"4A",X"49",X"48",X"47",X"46",X"46",X"45",X"44",X"44",X"43",X"43",X"42",X"41",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3C",X"3B",X"3B",X"3B",X"63",X"63",X"63",X"63",X"63",X"63",X"5E",X"5A",X"57",X"55",X"52",X"50",X"4F",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",X"46",X"46",X"45",X"44",X"44",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"3C",X"3B",X"63",X"63",X"63",X"63",X"63",X"63",X"5F",X"5B",X"58",X"55",X"53",X"51",X"4F",X"4E",X"4D",X"4B",X"4A",X"49",X"48",X"48",X"47",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3D",X"3C",X"3C",X"3C",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5C",X"59",X"56",X"54",X"52",X"50",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",X"47",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3D",X"3C",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5C",X"59",X"56",X"54",X"52",X"51",X"4F",X"4E",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"47",X"46",X"46",X"45",X"45",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3D",X"3D",X"3D",X"3D",X"63",X"63",X"63",X"63",X"63",X"63",X"61",X"5D",X"5A",X"57",X"55",X"53",X"51",X"50",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"48",X"47",X"46",X"46",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",X"3D",X"3D",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"5E",X"5A",X"58",X"55",X"53",X"52",X"50",X"4F",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"47",X"47",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"3E",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"5E",X"5B",X"58",X"56",X"54",X"52",X"51",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"48",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3F",X"3E",X"3E",X"3E",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"5F",X"5B",X"59",X"56",X"54",X"53",X"51",X"50",X"4E",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3F",X"3E",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"5F",X"5C",X"59",X"57",X"55",X"53",X"52",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"3F",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5C",X"5A",X"57",X"55",X"54",X"52",X"51",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"48",X"47",X"47",X"46",X"45",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"41",X"41",X"41",X"41",X"40",X"40",X"40",X"3F",X"3F",X"3F",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5D",X"5A",X"58",X"56",X"54",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"40",X"3F",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"61",X"5D",X"5B",X"58",X"56",X"54",X"53",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"40",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"61",X"5E",X"5B",X"59",X"57",X"55",X"53",X"52",X"51",X"4F",X"4E",X"4D",X"4C",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"40",X"40",X"40",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"5E",X"5C",X"59",X"57",X"55",X"54",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"41",X"40",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"5F",X"5C",X"5A",X"57",X"56",X"54",X"53",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"41",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"5F",X"5C",X"5A",X"58",X"56",X"54",X"53",X"52",X"51",X"4F",X"4E",X"4E",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"41",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5D",X"5A",X"58",X"56",X"55",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4C",X"4B",X"4A",X"4A",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"41",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5D",X"5B",X"59",X"57",X"55",X"54",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4D",X"4C",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"42",X"41",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"60",X"5E",X"5B",X"59",X"57",X"56",X"54",X"53",X"52",X"50",X"4F",X"4F",X"4E",X"4D",X"4C",X"4B",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"42",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"61",X"5E",X"5C",X"59",X"58",X"56",X"54",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4C",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"42",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"61",X"5E",X"5C",X"5A",X"58",X"56",X"55",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4E",X"4D",X"4C",X"4B",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"46",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43",X"42",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"63",X"62",X"5F",X"5C",X"5A",X"58",X"57",X"55",X"54",X"53",X"51",X"50",X"4F",X"4F",X"4E",X"4D",X"4C",X"4C",X"4B",X"4A",X"4A",X"49",X"49",X"48",X"48",X"47",X"47",X"47",X"46",X"46",X"46",X"45",X"45",X"45",X"44",X"44",X"44",X"43",X"43",X"43",X"43");
signal mult: ram_ir := (X"000",X"030",X"060",X"090",X"0C0",X"0F0",X"120",X"150",X"180",X"1B0",X"1E0",X"210",X"240",X"270",X"2A0",X"2D0",X"300",X"330",X"360",X"390",X"3C0",X"3F0",X"420",X"450",X"480",X"4B0",X"4E0",X"510",X"540",X"570",X"5A0",X"5D0",X"600",X"630",X"660",X"690",X"6C0",X"6F0",X"720",X"750",X"780",X"7B0",X"7E0",X"810",X"840",X"870",X"8A0",X"8D0");
signal shifted_sat : std_logic_vector(9 downto 0);
signal calibrated : integer := 0;
signal calibratedp30 : integer := 0;
signal diff : integer := 0;
signal modify : std_logic;
begin

--std_logic_vector(to_unsigned(ir, data_o'length));
	red_int <= "0000" & red_in(9 downto 4);
	ir_int <= "0000" & ir_in( 9 downto 4);
	red <= to_integer(unsigned(red_int));
	ir <= to_integer(unsigned(ir_int));
--	data_o <= std_logic_vector(to_unsigned(red_in,data_o'length)) when o_sel = '1' else std_logic_vector(to_unsigned(ir_in,data_o'length));
--   	data_o <= red_in when o_sel = '1' else ir_in;
	shifted_sat <= "00"&sat(ir + to_integer(unsigned(mult(red))));
	calibrated <= to_integer(unsigned(shifted_sat));
	calibratedp30 <= calibrated + 30;
	last_sat <= cur_sat;
	cur_sat <= std_logic_vector(to_unsigned(calibrated, data_o'length)) when calibrated > 69
		  else std_logic_vector(to_unsigned(calibratedp30, data_o'length));
	diff <= to_integer(unsigned(cur_sat)) - to_integer(unsigned(last_sat));
	modify <= '0' when diff > 10 
		else '0' when diff < -10
		else '1';
	sum_sat <= std_logic_vector(to_unsigned(to_integer(unsigned(cur_sat))+to_integer(unsigned(last_sat)),sum_sat'length)) when modify = '1' else last_sat;
	avg_sat <= "0" & sum_sat(9 downto 1);
	data_o <= cur_sat;end Behavioral;
